package wb_cov_pkg;

  import uvm_pkg::*;
  import wb_tlm_pkg::*;

  `include "uvm_macros.svh"
  `include "uvm_wb_queue.sv"
  `include "wb_cov.sv"

endpackage

