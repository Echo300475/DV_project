package wb_tlm_pkg;

  import uvm_pkg::*;

  `include "uvm_macros.svh"
  `include "wb_tlm.sv"

endpackage
