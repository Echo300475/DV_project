package wb_agent_pkg;
   
   import uvm_pkg::*;
   import wb_cfg_pkg::*;
   import wb_tlm_pkg::*;
   
   `include "uvm_macros.svh"
   `include "wb_master_driver_base.sv"
   `include "wb_master_driver.sv"
   `include "wb_slave_monitor.sv"
   `include "wb_agent.sv"
   
endpackage
