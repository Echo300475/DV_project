package wb_cfg_pkg;

  import uvm_pkg::*;

  `include "uvm_macros.svh"
  `include "wb_cfg.sv"

endpackage
