package wb_env_pkg;

  import uvm_pkg::*;
  import wb_agent_pkg::*;
  import wb_chk_pkg::*;
  import wb_cov_pkg::*;

  `include "uvm_macros.svh"
  `include "wb_env.svh"

endpackage