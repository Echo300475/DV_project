class wb_base_test extends uvm_test;

  `uvm_component_utils(wb_base_test)

  string my_name = "wb_base_test";

  typedef wb_env #(wb_tlm,wb_tlm) env_t;
  env_t env_h;
  wb_cfg wb_cfg_h;

  function new(string name, uvm_component parent);
    super.new(name,parent);
  endfunction

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    $display("-------------------------------------------------------------------------------------------------------------------------------------------");
    uvm_report_info(my_name, "base build phase");
    $display("-------------------------------------------------------------------------------------------------------------------------------------------");

    env_h = env_t::type_id::create("wb_env", this);
    $display("-------------------------------------------------------------------------------------------------------------------------------------------");
    `uvm_info(my_name,"env created",UVM_NONE)
    $display("-------------------------------------------------------------------------------------------------------------------------------------------");

    wb_cfg_h = wb_cfg::type_id::create("wb_cfg");
    $display("-------------------------------------------------------------------------------------------------------------------------------------------");
    `uvm_info(my_name,"wb_cfg created",UVM_NONE)
    $display("-------------------------------------------------------------------------------------------------------------------------------------------");

    uvm_config_db#(wb_cfg)::set(null,"*","WB_CFG",wb_cfg_h);
    $display("-------------------------------------------------------------------------------------------------------------------------------------------");
    `uvm_info(my_name,"wb_cfg is set into database",UVM_NONE)
    $display("-------------------------------------------------------------------------------------------------------------------------------------------");
  endfunction 

  function void start_of_simulation_phase(uvm_phase phase);
    $display("-------------------------------------------------------------------------------------------------------------------------------------------");
    uvm_report_info(my_name, "start of simulation");
    $display("-------------------------------------------------------------------------------------------------------------------------------------------");
  endfunction

endclass
