//***************************************************************************************************************
// Author: Van Le
// vanleatwork@yahoo.com
// Phone: VN: 0396221156, US: 5125841843
//***************************************************************************************************************
package spi_agent_pkg;
   
   import uvm_pkg::*;
   import spi_cfg_pkg::*;
   import spi_tlm_pkg::*;
   
   `include "uvm_macros.svh"
   //`include "spi_monitor.sv"
   `include "spi_driver_base.sv"
   `include "spi_driver.sv"
   `include "spi_agent.sv"

endpackage
