package wb_seq_pkg;

   import uvm_pkg::*;
   import wb_cfg_pkg::*;
   import wb_tlm_pkg::*;

   `include "uvm_macros.svh"
   `include "base_seq.sv"
   `include "rst_seq.sv"
   `include "wb_single_wr_rd.sv"
   `include "wb_block_wr_rd.sv"

endpackage
