package wb_chk_pkg;

  import uvm_pkg::*;
  import wb_tlm_pkg::*;
  import wb_cfg_pkg::*;

  `include "uvm_macros.svh"
  `include "sb.sv"

endpackage
